`timescale 1ns / 1ps

module tb;

   reg [7:0] sw;
   reg       clk;
   reg       btnS;
   reg       btnR;
   
   integer   i;
   
   /*AUTOWIRE*/
   // Beginning of automatic wires (for undeclared instantiated-module outputs)
   wire                 RsRx;                   // From model_uart0_ of model_uart.v
   wire                 RsTx;                   // From uut_ of nexys3.v
   wire [7:0]           led;                    // From uut_ of nexys3.v
   // End of automatics

   /* For reading */
   integer file;
   integer numlines;
   reg [7:0] mem [0:1024];
   integer j;
   integer reg1;
   integer reg2;
   integer reg3;
   integer pushed;
   
   initial
     begin
        //$shm_open  ("dump", , ,1);
        //$shm_probe (tb, "ASTF");

        clk = 0;
        btnR = 1;
        btnS = 0;
        btnR = 0;
		#100
		// Read in code
		
		file = $fopen("seq.code", "rb");
		
		$fscanf(file, "%b\n", numlines);
		$readmemb("seq.code", mem);
		
		j = 1;
		repeat (numlines) begin
			if (mem[j][7] == 0 && mem[j][6] == 0) begin
				reg1 = 2* mem[j][5] + mem[j][4];
				pushed = 8 * mem[j][3] + 4 * mem[j][2] + 2 * mem[j][1] + mem[j][0];
				tskRunPUSH(reg1, pushed);
				
			end
			
			else if (mem[j][7] == 0 && mem[j][6] == 1) begin
				reg1 = 2* mem[j][5] + mem[j][4];
				reg2 = 2* mem[j][3] + mem[j][2];
				reg3 = 2* mem[j][1] + mem[j][0];
				tskRunADD(reg1, reg2, reg3);
			end
			
			else if (mem[j][7] == 1 && mem[j][6] == 0) begin
				
				reg1 = 2* mem[j][5] + mem[j][4];
				reg2 = 2* mem[j][3] + mem[j][2];
				reg3 = 2* mem[j][1] + mem[j][0];
				tskRunMULT(reg1, reg2, reg3);
			end
			
			
			else if (mem[j][7] == 1 && mem[j][6] == 1) begin
				
				reg1 = 2* mem[j][5] + mem[j][4];
				tskRunSEND(reg1);
				$display("SENDING");
			end
			j = j + 1;
		end
		
		/*
        tskRunPUSH(0,4);
        tskRunPUSH(0,0);
        tskRunPUSH(1,3);
        tskRunMULT(0,1,2);
        tskRunADD(2,0,3);
        tskRunSEND(0);
        tskRunSEND(1);
        tskRunSEND(2);
        tskRunSEND(3); */
        
        #1500000000;     
		$display("Done");
        $finish;
     end

   always #5 clk = ~clk;
   
   model_uart model_uart0_ (// Outputs
                            .TX                  (RsRx),
                            // Inputs
                            .RX                  (RsTx)
                            /*AUTOINST*/);

   defparam model_uart0_.name = "UART0";
   defparam model_uart0_.baud = 1000000;
   
   
   nexys3 uut_ (/*AUTOINST*/
                // Outputs
                .RsTx                   (RsTx),
                .led                    (led[7:0]),
                // Inputs
                .RsRx                   (RsRx),
                .sw                     (sw[7:0]),
                .btnS                   (btnS),
                .btnR                   (btnR),
                .clk                    (clk));

   task tskRunInst;
      input [7:0] inst;
      begin
         $display ("%d ... Running instruction %08b", $stime, inst);
         sw = inst;
         #1500000 btnS = 1;
         #3000000 btnS = 0;
      end
   endtask //

   task tskRunPUSH;
      input [1:0] ra;
      input [3:0] immd;
      reg [7:0]   inst;
      begin
         inst = {2'b00, ra[1:0], immd[3:0]};
         tskRunInst(inst);
      end
   endtask //

   task tskRunSEND;
      input [1:0] ra;
      reg [7:0]   inst;
      begin
         inst = {2'b11, ra[1:0], 4'h0};
         tskRunInst(inst);
      end
   endtask //

   task tskRunADD;
      input [1:0] ra;
      input [1:0] rb;
      input [1:0] rc;
      reg [7:0]   inst;
      begin
         inst = {2'b01, ra[1:0], rb[1:0], rc[1:0]};
         tskRunInst(inst);
      end
   endtask //

   task tskRunMULT;
      input [1:0] ra;
      input [1:0] rb;
      input [1:0] rc;
      reg [7:0]   inst;
      begin
         inst = {2'b10, ra[1:0], rb[1:0], rc[1:0]};
         tskRunInst(inst);
      end
   endtask //

   always @ (posedge clk)
     if (uut_.inst_vld)
       $display("%d ... instruction %08b executed", $stime, uut_.inst_wd);

   always @ (led)
     $display("%d ... led output changed to %08b", $stime, led);
   
endmodule // tb
// Local Variables:
// verilog-library-flags:("-y ../src/")
// End:
